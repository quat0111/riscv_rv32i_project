
`timescale 1ns/1ps

module tb_Control_Logic;

    // Inputs
    logic [31:0] instr;
    logic        BrEq;
    logic        BrLT;

    // Outputs
    logic        PCSel;
    logic [2:0]  ImmSel;
    logic        RegWEn;
    logic        BrUn;
    logic        BSel;
    logic        ASel;
    logic [3:0]  ALUSel;
    logic        MemRW;
    logic [1:0]  WBSel;

    // DUT
    Control_Logic ctrl (
        .instr(instr),
        .PCSel(PCSel),
        .BrEq(BrEq),
        .BrLT(BrLT),
        .RegWEn(RegWEn),
        .BrUn(BrUn),
        .Bsel(BSel),
        .Asel(ASel),
        .MemRW(MemRW),
        .ImmSel(ImmSel),
        .ALUSel(ALUSel),
        .WBSel(WBSel)
    );

    initial begin
        BrEq = 0;
        BrLT = 0;

        // ============================================================
        // R-TYPE (ADD x1, x2, x3)
        // opcode 0x33, funct3=0, funct7=0  → ADD
        // ============================================================
        instr = 32'h003100B3;   // ADD x1, x2, x3
        #10;

        // ============================================================
        // I-TYPE (ADDI x1, x2, 5)
        // opcode 0x13
        // ============================================================
        instr = 32'h00510093;   // ADDI x1, x2, 5
        #10;

        // ============================================================
        // LOAD (LW x1, 4(x2))
        // opcode 0x03, funct3 = 010
        // ============================================================
        instr = 32'h00412083;   // LW x1, 4(x2)
        #10;

        // ============================================================
        // STORE (SW x1, 4(x2))
        // opcode 0x23
        // ============================================================
        instr = 32'h00112223;   // SW x1, 4(x2)
        #10;

        // ============================================================
        // BRANCH: BEQ x1, x2, offset
        // ============================================================
        BrEq = 1;
        instr = 32'h00208863;   // BEQ (taken)
        #10;
        BrEq = 0;               // BEQ (not taken)
        #10;

        // ============================================================
        // JAL (jump and link)
        // ============================================================
        instr = 32'h00c000ef;   // JAL x1, 12
        #10;

        // ============================================================
        // JALR (jump register)
        // ============================================================
        instr = 32'h004100E7;   // JALR x1, 4(x2)
        #10;

        // ============================================================
        // LUI x1, imm
        // ============================================================
        instr = 32'h000010B7;   // LUI x1, 0x1
        #10;

        // ============================================================
        // AUIPC x1, imm
        // ============================================================
        instr = 32'h00001097;   // AUIPC x1, 0x1
        #10;

        $finish;
    end

endmodule
